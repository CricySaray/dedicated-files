//-----------------------------------------------------------------------------
// Company: QUST
// Engineer: 宋安瑞
//
// Create Date: 2022年9月14日15:53:20
// Design Name: 6_64decoder
// Module Name: design file
// Target Device: any
// Tool versions: any
// Description:
// 				
// Dependencies: 
// 				
// Revision:
// 				
// Additional Comments:
// 
//-----------------------------------------------------------------------------

`timescale 1ns/1ns

module decoder6_64_sar(in, out);
	input [0:5] in;
	output [0:63] out;
	reg [0:63] out;

	always @(in) 
		begin 
			case (in)
				6'b000_000 : out=64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001;
				6'b000_001 : out=64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010;
				6'b000_010 : out=64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100;
				6'b000_011 : out=64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000;
				6'b000_100 : out=64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00010000;
				6'b000_101 : out=64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00100000;
				6'b000_110 : out=64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_01000000;
				6'b000_111 : out=64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000;

				6'b001_000 : out=64'b00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000;
				6'b001_001 : out=64'b00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000;
				6'b001_010 : out=64'b00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000;
				6'b001_011 : out=64'b00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000;
				6'b001_100 : out=64'b00000000_00000000_00000000_00000000_00000000_00000000_00010000_00000000;
				6'b001_101 : out=64'b00000000_00000000_00000000_00000000_00000000_00000000_00100000_00000000;
				6'b001_110 : out=64'b00000000_00000000_00000000_00000000_00000000_00000000_01000000_00000000;
				6'b001_111 : out=64'b00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000;

				6'b010_000 : out=64'b00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000;
				6'b010_001 : out=64'b00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000;
				6'b010_010 : out=64'b00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000;
				6'b010_011 : out=64'b00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000;
				6'b010_100 : out=64'b00000000_00000000_00000000_00000000_00000000_00010000_00000000_00000000;
				6'b010_101 : out=64'b00000000_00000000_00000000_00000000_00000000_00100000_00000000_00000000;
				6'b010_110 : out=64'b00000000_00000000_00000000_00000000_00000000_01000000_00000000_00000000;
				6'b010_111 : out=64'b00000000_00000000_00000000_00000000_00000000_10000000_00000000_00000000;

				6'b011_000 : out=64'b00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000;
				6'b011_001 : out=64'b00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000;
				6'b011_010 : out=64'b00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000;
				6'b011_011 : out=64'b00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000;
				6'b011_100 : out=64'b00000000_00000000_00000000_00000000_00010000_00000000_00000000_00000000;
				6'b011_101 : out=64'b00000000_00000000_00000000_00000000_00100000_00000000_00000000_00000000;
				6'b011_110 : out=64'b00000000_00000000_00000000_00000000_01000000_00000000_00000000_00000000;
				6'b011_111 : out=64'b00000000_00000000_00000000_00000000_10000000_00000000_00000000_00000000;

				6'b100_000 : out=64'b00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000;
				6'b100_001 : out=64'b00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000;
				6'b100_010 : out=64'b00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000;
				6'b100_011 : out=64'b00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000;
				6'b100_100 : out=64'b00000000_00000000_00000000_00010000_00000000_00000000_00000000_00000000;
				6'b100_101 : out=64'b00000000_00000000_00000000_00100000_00000000_00000000_00000000_00000000;
				6'b100_110 : out=64'b00000000_00000000_00000000_01000000_00000000_00000000_00000000_00000000;
				6'b100_111 : out=64'b00000000_00000000_00000000_10000000_00000000_00000000_00000000_00000000;

				6'b101_000 : out=64'b00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000;
				6'b101_001 : out=64'b00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000;
				6'b101_010 : out=64'b00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000;
				6'b101_011 : out=64'b00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000;
				6'b101_100 : out=64'b00000000_00000000_00010000_00000000_00000000_00000000_00000000_00000000;
				6'b101_101 : out=64'b00000000_00000000_00100000_00000000_00000000_00000000_00000000_00000000;
				6'b101_110 : out=64'b00000000_00000000_01000000_00000000_00000000_00000000_00000000_00000000;
				6'b101_111 : out=64'b00000000_00000000_10000000_00000000_00000000_00000000_00000000_00000000;

				6'b110_000 : out=64'b00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000;
				6'b110_001 : out=64'b00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000;
				6'b110_010 : out=64'b00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000;
				6'b110_011 : out=64'b00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000;
				6'b110_100 : out=64'b00000000_00010000_00000000_00000000_00000000_00000000_00000000_00000000;
				6'b110_101 : out=64'b00000000_00100000_00000000_00000000_00000000_00000000_00000000_00000000;
				6'b110_110 : out=64'b00000000_01000000_00000000_00000000_00000000_00000000_00000000_00000000;
				6'b110_111 : out=64'b00000000_10000000_00000000_00000000_00000000_00000000_00000000_00000000;

				6'b111_000 : out=64'b00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
				6'b111_001 : out=64'b00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
				6'b111_010 : out=64'b00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
				6'b111_011 : out=64'b00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
				6'b111_100 : out=64'b00010000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
				6'b111_101 : out=64'b00100000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
				6'b111_110 : out=64'b01000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
				6'b111_111 : out=64'b10000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;

				
				default: out=64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
			endcase
		end
endmodule 
		