module decoder(decoderout,waddr);
output[31:0] decoderout;
input[4:0] waddr;

reg [31:0] decoderout;

always @ (waddr)
case(waddr)
5'd0: decoderout=32'b0000_0000_0000_0000_0000_0000_0000_0001;
5'd1: decoderout=32'b0000_0000_0000_0000_0000_0000_0000_0010;
5'd2: decoderout=32'b0000_0000_0000_0000_0000_0000_0000_0100;
5'd3: decoderout=32'b0000_0000_0000_0000_0000_0000_0000_1000;
5'd4: decoderout=32'b0000_0000_0000_0000_0000_0000_0001_0000;
5'd5: decoderout=32'b0000_0000_0000_0000_0000_0000_0010_0000;
5'd6: decoderout=32'b0000_0000_0000_0000_0000_0000_0100_0000;
5'd7: decoderout=32'b0000_0000_0000_0000_0000_0000_1000_0000;
5'd8: decoderout=32'b0000_0000_0000_0000_0000_0001_0000_0000;
5'd9: decoderout=32'b0000_0000_0000_0000_0000_0010_0000_0000;
5'd10: decoderout=32'b0000_0000_0000_0000_0000_0100_0000_0000;
5'd11: decoderout=32'b0000_0000_0000_0000_0000_1000_0000_0000;
5'd12: decoderout=32'b0000_0000_0000_0000_0001_0000_0000_0000;
5'd13: decoderout=32'b0000_0000_0000_0000_0010_0000_0000_0000;
5'd14: decoderout=32'b0000_0000_0000_0000_0100_0000_0000_0000;
5'd15: decoderout=32'b0000_0000_0000_0000_1000_0000_0000_0000;
5'd16: decoderout=32'b0000_0000_0000_0001_0000_0000_0000_0000;
5'd17: decoderout=32'b0000_0000_0000_0010_0000_0000_0000_0000;
5'd18: decoderout=32'b0000_0000_0000_0100_0000_0000_0000_0000;
5'd19: decoderout=32'b0000_0000_0000_1000_0000_0000_0000_0000;
5'd20: decoderout=32'b0000_0000_0001_0000_0000_0000_0000_0000;
5'd21: decoderout=32'b0000_0000_0010_0000_0000_0000_0000_0000;
5'd22: decoderout=32'b0000_0000_0100_0000_0000_0000_0000_0000;
5'd23: decoderout=32'b0000_0000_1000_0000_0000_0000_0000_0000;
5'd24: decoderout=32'b0000_0001_0000_0000_0000_0000_0000_0000;
5'd25: decoderout=32'b0000_0010_0000_0000_0000_0000_0000_0000;
5'd26: decoderout=32'b0000_0100_0000_0000_0000_0000_0000_0000;
5'd27: decoderout=32'b0000_1000_0000_0000_0000_0000_0000_0000;
5'd28: decoderout=32'b0001_0000_0000_0000_0000_0000_0000_0000;
5'd29: decoderout=32'b0010_0000_0000_0000_0000_0000_0000_0000;
5'd30: decoderout=32'b0100_0000_0000_0000_0000_0000_0000_0000;
5'd31: decoderout=32'b1000_0000_0000_0000_0000_0000_0000_0000;
endcase
endmodule